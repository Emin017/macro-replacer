module NEW_MACRO(
  input CLK,
  input WEN,
  input [3:0] D,
  output [3:0] Q
);
endmodule
