module NEW_MACRO(input X, input Y); endmodule
