module top;
  OLD_MACRO u_inst (.A(a), .B(b));
endmodule
